module clock_divider(
	input clock,
	output imem_clock, 
	output dmem_clock, 
	output processor_clock, 
	output regfile_clock
);



endmodule
